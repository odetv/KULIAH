CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1918 1029
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
58
13 Logic Switch~
5 146 99 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -16 7 -8
2 D1
-6 -26 8 -18
9 SERIAL IN
-31 -36 32 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90023e-315 0
0
13 Logic Switch~
5 69 98 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-7 -15 7 -7
2 V4
-7 -25 7 -17
5 CLOCK
-17 -36 18 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90023e-315 5.26354e-315
0
9 Inverter~
13 217 1521 0 2 22
0 7 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U20E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 16 0
1 U
3124 0 0
2
5.90023e-315 5.45782e-315
0
10 2-In NAND~
219 296 1417 0 3 22
0 7 6 12
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U23D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
3421 0 0
2
5.90023e-315 5.45523e-315
0
10 2-In NAND~
219 295 1512 0 3 22
0 6 9 11
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
8157 0 0
2
5.90023e-315 5.45264e-315
0
10 2-In NAND~
219 438 1503 0 3 22
0 2 11 10
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 20 0
1 U
5572 0 0
2
5.90023e-315 5.45005e-315
0
10 2-In NAND~
219 437 1426 0 3 22
0 12 10 2
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 20 0
1 U
8901 0 0
2
5.90023e-315 5.44746e-315
0
14 Logic Display~
6 1051 99 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.90023e-315 5.44487e-315
0
14 Logic Display~
6 561 1481 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.90023e-315 5.44228e-315
0
9 Inverter~
13 215 1333 0 2 22
0 5 13
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U20F
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 16 0
1 U
972 0 0
2
5.90023e-315 5.43969e-315
0
10 2-In NAND~
219 294 1229 0 3 22
0 5 6 16
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 20 0
1 U
3472 0 0
2
5.90023e-315 5.4371e-315
0
10 2-In NAND~
219 293 1324 0 3 22
0 6 13 15
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
9998 0 0
2
5.90023e-315 5.43451e-315
0
10 2-In NAND~
219 436 1315 0 3 22
0 7 15 14
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
3536 0 0
2
5.90023e-315 5.43192e-315
0
10 2-In NAND~
219 435 1238 0 3 22
0 16 14 7
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 21 0
1 U
4597 0 0
2
5.90023e-315 5.42933e-315
0
14 Logic Display~
6 1003 98 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.90023e-315 5.42414e-315
0
14 Logic Display~
6 559 1293 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90023e-315 5.41896e-315
0
14 Logic Display~
6 557 1107 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90023e-315 5.41378e-315
0
14 Logic Display~
6 954 97 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.90023e-315 5.4086e-315
0
10 2-In NAND~
219 433 1052 0 3 22
0 20 18 5
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 21 0
1 U
317 0 0
2
5.90023e-315 5.40342e-315
0
10 2-In NAND~
219 434 1129 0 3 22
0 5 19 18
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
3108 0 0
2
5.90023e-315 5.39824e-315
0
10 2-In NAND~
219 291 1138 0 3 22
0 6 17 19
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 22 0
1 U
4299 0 0
2
5.90023e-315 5.39306e-315
0
10 2-In NAND~
219 292 1043 0 3 22
0 8 6 20
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 22 0
1 U
9672 0 0
2
5.90023e-315 5.38788e-315
0
9 Inverter~
13 213 1147 0 2 22
0 8 17
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 23 0
1 U
7876 0 0
2
5.90023e-315 5.37752e-315
0
9 Inverter~
13 212 955 0 2 22
0 3 21
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 23 0
1 U
6369 0 0
2
5.90023e-315 5.36716e-315
0
10 2-In NAND~
219 291 851 0 3 22
0 3 6 24
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 22 0
1 U
9172 0 0
2
5.90023e-315 5.3568e-315
0
10 2-In NAND~
219 290 946 0 3 22
0 6 21 23
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 24 0
1 U
7100 0 0
2
5.90023e-315 5.34643e-315
0
10 2-In NAND~
219 433 937 0 3 22
0 8 23 22
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 24 0
1 U
3820 0 0
2
5.90023e-315 5.32571e-315
0
10 2-In NAND~
219 432 860 0 3 22
0 24 22 8
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 24 0
1 U
7678 0 0
2
5.90023e-315 5.30499e-315
0
14 Logic Display~
6 907 95 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90023e-315 5.26354e-315
0
14 Logic Display~
6 556 915 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
5.90023e-315 0
0
9 Inverter~
13 212 778 0 2 22
0 25 27
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U20D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 16 0
1 U
3409 0 0
2
5.90023e-315 5.30499e-315
0
10 2-In NAND~
219 291 674 0 3 22
0 25 6 30
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U23C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
3951 0 0
2
5.90023e-315 5.32571e-315
0
10 2-In NAND~
219 290 769 0 3 22
0 6 27 29
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U23B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 19 0
1 U
8885 0 0
2
5.90023e-315 5.34643e-315
0
10 2-In NAND~
219 433 760 0 3 22
0 3 29 28
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U23A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 19 0
1 U
3780 0 0
2
5.90023e-315 5.3568e-315
0
10 2-In NAND~
219 432 683 0 3 22
0 30 28 3
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U22D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
9265 0 0
2
5.90023e-315 5.36716e-315
0
14 Logic Display~
6 858 95 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L28
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
5.90023e-315 5.37752e-315
0
14 Logic Display~
6 556 738 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L27
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
5.90023e-315 5.38788e-315
0
9 Inverter~
13 210 590 0 2 22
0 4 31
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U20C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 16 0
1 U
9968 0 0
2
5.90023e-315 5.39306e-315
0
10 2-In NAND~
219 289 486 0 3 22
0 4 6 34
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U22C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
9281 0 0
2
5.90023e-315 5.39824e-315
0
10 2-In NAND~
219 288 581 0 3 22
0 6 31 33
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U22B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
8464 0 0
2
5.90023e-315 5.40342e-315
0
10 2-In NAND~
219 431 572 0 3 22
0 25 33 32
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U22A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
7168 0 0
2
5.90023e-315 5.4086e-315
0
10 2-In NAND~
219 430 495 0 3 22
0 34 32 25
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U21D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
3171 0 0
2
5.90023e-315 5.41378e-315
0
14 Logic Display~
6 805 95 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.90023e-315 5.41896e-315
0
14 Logic Display~
6 554 550 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6435 0 0
2
5.90023e-315 5.42414e-315
0
14 Logic Display~
6 552 364 0 1 2
10 36
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
5.90023e-315 5.42933e-315
0
14 Logic Display~
6 750 97 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
5.90023e-315 5.43192e-315
0
10 2-In NAND~
219 428 309 0 3 22
0 38 36 4
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U21C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
5305 0 0
2
5.90023e-315 5.43451e-315
0
10 2-In NAND~
219 429 386 0 3 22
0 4 37 36
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U21B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
34 0 0
2
5.90023e-315 5.4371e-315
0
10 2-In NAND~
219 286 395 0 3 22
0 6 35 37
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U21A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
969 0 0
2
5.90023e-315 5.43969e-315
0
10 2-In NAND~
219 287 300 0 3 22
0 26 6 38
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
8402 0 0
2
5.90023e-315 5.44228e-315
0
9 Inverter~
13 208 404 0 2 22
0 26 35
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U20B
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 16 0
1 U
3751 0 0
2
5.90023e-315 5.44487e-315
0
9 Inverter~
13 207 212 0 2 22
0 39 40
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U20A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 16 0
1 U
4292 0 0
2
5.90023e-315 5.44746e-315
0
10 2-In NAND~
219 286 108 0 3 22
0 39 6 43
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
6118 0 0
2
5.90023e-315 5.45005e-315
0
10 2-In NAND~
219 285 203 0 3 22
0 6 40 42
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
34 0 0
2
5.90023e-315 5.45264e-315
0
10 2-In NAND~
219 428 194 0 3 22
0 26 42 41
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
6357 0 0
2
5.90023e-315 5.45523e-315
0
10 2-In NAND~
219 427 117 0 3 22
0 43 41 26
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
319 0 0
2
5.90023e-315 5.45782e-315
0
14 Logic Display~
6 697 98 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
5.90023e-315 5.46041e-315
0
14 Logic Display~
6 551 172 0 1 2
10 41
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
5.90023e-315 5.463e-315
0
88
0 1 2 0 0 8192 0 0 6 17 0 5
497 1426
497 1468
403 1468
403 1494
414 1494
1 0 3 0 0 12288 0 34 0 0 58 5
409 751
399 751
399 726
492 726
492 683
0 0 4 0 0 8320 0 0 0 76 61 4
594 309
594 435
185 435
185 477
0 0 5 0 0 8192 0 0 0 35 20 4
597 1052
597 1180
190 1180
190 1220
0 0 6 0 0 8192 0 0 0 19 6 3
255 1463
83 1463
83 1277
0 0 6 0 0 8192 0 0 0 28 7 3
253 1277
83 1277
83 1090
0 0 6 0 0 8192 0 0 0 37 8 3
251 1090
83 1090
83 899
0 0 6 0 0 0 0 0 0 46 48 3
250 899
83 899
83 719
1 0 3 0 0 0 0 25 0 0 38 2
267 842
187 842
0 0 7 0 0 8192 0 0 0 26 12 4
599 1238
599 1368
192 1368
192 1408
0 0 8 0 0 8192 0 0 0 44 29 4
598 860
598 1003
188 1003
188 1036
1 1 7 0 0 0 0 3 4 0 0 4
202 1521
192 1521
192 1408
272 1408
2 2 9 0 0 4224 0 5 3 0 0 2
271 1521
238 1521
2 0 10 0 0 12288 0 7 0 0 15 5
413 1435
404 1435
404 1459
483 1459
483 1503
3 1 10 0 0 4224 0 6 9 0 0 3
465 1503
561 1503
561 1499
3 2 11 0 0 4224 0 5 6 0 0 2
322 1512
414 1512
3 1 2 0 0 8320 0 7 8 0 0 3
464 1426
1051 1426
1051 117
3 1 12 0 0 4224 0 4 7 0 0 2
323 1417
413 1417
1 2 6 0 0 0 0 5 4 0 0 4
271 1503
255 1503
255 1426
272 1426
1 1 5 0 0 0 0 10 11 0 0 4
200 1333
190 1333
190 1220
270 1220
2 2 13 0 0 4224 0 12 10 0 0 2
269 1333
236 1333
2 0 14 0 0 12288 0 14 0 0 23 5
411 1247
402 1247
402 1271
481 1271
481 1315
3 1 14 0 0 4224 0 13 16 0 0 3
463 1315
559 1315
559 1311
3 2 15 0 0 4224 0 12 13 0 0 2
320 1324
412 1324
1 0 7 0 0 0 0 13 0 0 26 5
412 1306
402 1306
402 1281
494 1281
494 1238
3 1 7 0 0 8320 0 14 15 0 0 3
462 1238
1003 1238
1003 116
3 1 16 0 0 4224 0 11 14 0 0 2
321 1229
411 1229
1 2 6 0 0 0 0 12 11 0 0 4
269 1315
253 1315
253 1238
270 1238
1 1 8 0 0 0 0 23 22 0 0 4
198 1147
188 1147
188 1034
268 1034
2 2 17 0 0 4224 0 21 23 0 0 2
267 1147
234 1147
2 0 18 0 0 12288 0 19 0 0 32 5
409 1061
400 1061
400 1085
479 1085
479 1129
3 1 18 0 0 4224 0 20 17 0 0 3
461 1129
557 1129
557 1125
3 2 19 0 0 4224 0 21 20 0 0 2
318 1138
410 1138
1 0 5 0 0 0 0 20 0 0 35 5
410 1120
400 1120
400 1095
492 1095
492 1052
3 1 5 0 0 8320 0 19 18 0 0 3
460 1052
954 1052
954 115
3 1 20 0 0 4224 0 22 19 0 0 2
319 1043
409 1043
1 2 6 0 0 0 0 21 22 0 0 4
267 1129
251 1129
251 1052
268 1052
1 0 3 0 0 12288 0 24 0 0 58 5
197 955
187 955
187 814
600 814
600 683
2 2 21 0 0 4224 0 26 24 0 0 2
266 955
233 955
2 0 22 0 0 12288 0 28 0 0 41 5
408 869
399 869
399 893
478 893
478 937
3 1 22 0 0 4224 0 27 30 0 0 3
460 937
556 937
556 933
3 2 23 0 0 4224 0 26 27 0 0 2
317 946
409 946
1 0 8 0 0 0 0 27 0 0 44 5
409 928
399 928
399 903
491 903
491 860
3 1 8 0 0 8320 0 28 29 0 0 3
459 860
907 860
907 113
3 1 24 0 0 4224 0 25 28 0 0 2
318 851
408 851
1 2 6 0 0 0 0 26 25 0 0 4
266 937
250 937
250 860
267 860
0 0 25 0 0 8320 0 0 0 67 53 4
598 495
598 625
187 625
187 665
0 0 6 0 0 0 0 0 0 60 50 3
250 719
83 719
83 531
1 0 6 0 0 0 0 2 0 0 87 4
81 98
83 98
83 154
245 154
0 0 6 0 0 0 0 0 0 69 51 3
248 531
83 531
83 347
0 0 6 0 0 4224 0 0 0 49 78 3
83 154
83 347
246 347
0 0 26 0 0 8320 0 0 0 85 70 4
593 117
593 260
183 260
183 293
1 1 25 0 0 0 0 31 32 0 0 4
197 778
187 778
187 665
267 665
2 2 27 0 0 4224 0 33 31 0 0 2
266 778
233 778
2 0 28 0 0 12288 0 35 0 0 56 5
408 692
399 692
399 716
478 716
478 760
3 1 28 0 0 4224 0 34 37 0 0 3
460 760
556 760
556 756
3 2 29 0 0 4224 0 33 34 0 0 2
317 769
409 769
3 1 3 0 0 8320 0 35 36 0 0 3
459 683
858 683
858 113
3 1 30 0 0 4224 0 32 35 0 0 2
318 674
408 674
1 2 6 0 0 0 0 33 32 0 0 4
266 760
250 760
250 683
267 683
1 1 4 0 0 0 0 38 39 0 0 4
195 590
185 590
185 477
265 477
2 2 31 0 0 4224 0 40 38 0 0 2
264 590
231 590
2 0 32 0 0 12288 0 42 0 0 64 5
406 504
397 504
397 528
476 528
476 572
3 1 32 0 0 4224 0 41 44 0 0 3
458 572
554 572
554 568
3 2 33 0 0 4224 0 40 41 0 0 2
315 581
407 581
1 0 25 0 0 0 0 41 0 0 67 5
407 563
397 563
397 538
489 538
489 495
3 1 25 0 0 0 0 42 43 0 0 3
457 495
805 495
805 113
3 1 34 0 0 4224 0 39 42 0 0 2
316 486
406 486
1 2 6 0 0 0 0 40 39 0 0 4
264 572
248 572
248 495
265 495
1 1 26 0 0 0 0 51 50 0 0 4
193 404
183 404
183 291
263 291
2 2 35 0 0 4224 0 49 51 0 0 2
262 404
229 404
2 0 36 0 0 12288 0 47 0 0 73 5
404 318
395 318
395 342
474 342
474 386
3 1 36 0 0 4224 0 48 45 0 0 3
456 386
552 386
552 382
3 2 37 0 0 4224 0 49 48 0 0 2
313 395
405 395
1 0 4 0 0 0 0 48 0 0 76 5
405 377
395 377
395 352
487 352
487 309
3 1 4 0 0 0 0 47 46 0 0 3
455 309
750 309
750 115
3 1 38 0 0 4224 0 50 47 0 0 2
314 300
404 300
1 2 6 0 0 0 0 49 50 0 0 4
262 386
246 386
246 309
263 309
1 0 39 0 0 8320 0 52 0 0 88 3
192 212
182 212
182 99
2 2 40 0 0 4224 0 54 52 0 0 2
261 212
228 212
2 0 41 0 0 12288 0 56 0 0 82 5
403 126
394 126
394 150
473 150
473 194
3 1 41 0 0 4224 0 55 58 0 0 3
455 194
551 194
551 190
3 2 42 0 0 4224 0 54 55 0 0 2
312 203
404 203
1 0 26 0 0 0 0 55 0 0 85 5
404 185
394 185
394 160
486 160
486 117
3 1 26 0 0 0 0 56 57 0 0 3
454 117
697 117
697 116
3 1 43 0 0 4224 0 53 56 0 0 2
313 108
403 108
1 2 6 0 0 0 0 54 53 0 0 4
261 194
245 194
245 117
262 117
1 1 39 0 0 0 0 1 53 0 0 2
158 99
262 99
26
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
836 18 933 42
844 26 924 42
10 SERIAL OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
554 162 585 184
561 169 577 185
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
552 88 575 110
559 95 567 111
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
553 280 576 302
560 287 568 303
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
555 354 586 376
562 361 578 377
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
557 540 588 562
564 547 580 563
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
555 466 578 488
562 473 570 489
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
559 728 590 750
566 735 582 751
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
557 654 580 676
564 661 572 677
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
682 42 713 64
689 50 705 66
2 Q1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
735 43 768 65
743 50 759 66
2 Q2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
790 43 821 65
797 50 813 66
2 Q3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
843 44 876 66
851 51 867 67
2 Q4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
559 905 590 927
566 912 582 928
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
557 831 580 853
564 838 572 854
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
558 1023 581 1045
565 1030 573 1046
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
560 1097 591 1119
567 1104 583 1120
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
562 1283 593 1305
569 1290 585 1306
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
560 1209 583 1231
567 1216 575 1232
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
564 1471 595 1493
571 1478 587 1494
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
562 1397 585 1419
569 1404 577 1420
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
893 42 923 66
901 51 914 67
2 Q5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
942 47 967 71
946 51 962 67
2 Q6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
991 46 1016 70
995 50 1011 66
2 Q7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1039 47 1064 71
1043 51 1059 67
2 Q8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 43
41 20 347 44
50 28 337 44
43 RANGKAIAN REGISTER SISO 8 BIT (D FLIP-FLOP)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
