CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1918 1029
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
98
13 Logic Switch~
5 81 111 0 1 11
0 2
0
0 0 21856 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
5 CLOCK
-17 -36 18 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44633.6 0
0
13 Logic Switch~
5 206 111 0 10 11
0 83 0 0 0 0 0 0 0 0
1
0
0 0 21856 0
2 5V
-6 -16 8 -8
2 V7
-6 -26 8 -18
9 SERIAL IN
-31 -36 32 -28
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
44633.6 1
0
14 Logic Display~
6 890 1015 0 1 2
10 35
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
44633.6 2
0
9 Inverter~
13 432 1095 0 2 22
0 2 38
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U12E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3421 0 0
2
44633.6 3
0
10 2-In NAND~
219 656 957 0 3 22
0 38 41 37
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
8157 0 0
2
44633.6 4
0
10 2-In NAND~
219 656 1052 0 3 22
0 39 38 36
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5572 0 0
2
44633.6 5
0
10 2-In NAND~
219 800 1043 0 3 22
0 7 36 35
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
8901 0 0
2
44633.6 6
0
10 2-In NAND~
219 800 966 0 3 22
0 37 35 7
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
7361 0 0
2
44633.6 7
0
10 2-In NAND~
219 509 966 0 3 22
0 42 39 41
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
4747 0 0
2
44633.6 8
0
10 2-In NAND~
219 510 1043 0 3 22
0 41 40 39
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
972 0 0
2
44633.6 9
0
10 2-In NAND~
219 367 1052 0 3 22
0 2 43 40
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3472 0 0
2
44633.6 10
0
10 2-In NAND~
219 368 957 0 3 22
0 3 2 42
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
9998 0 0
2
44633.6 11
0
9 Inverter~
13 279 998 0 2 22
0 3 43
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U12F
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3536 0 0
2
44633.6 12
0
9 Inverter~
13 279 1209 0 2 22
0 7 34
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U6A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 15 0
1 U
4597 0 0
2
44633.6 13
0
10 2-In NAND~
219 368 1168 0 3 22
0 7 2 33
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
3835 0 0
2
44633.6 14
0
10 2-In NAND~
219 367 1263 0 3 22
0 2 34 31
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
3670 0 0
2
44633.6 15
0
10 2-In NAND~
219 510 1254 0 3 22
0 32 31 30
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
5616 0 0
2
44633.6 16
0
10 2-In NAND~
219 509 1177 0 3 22
0 33 30 32
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
9323 0 0
2
44633.6 17
0
10 2-In NAND~
219 800 1177 0 3 22
0 28 26 6
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
317 0 0
2
44633.6 18
0
10 2-In NAND~
219 800 1254 0 3 22
0 6 27 26
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U7D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
3108 0 0
2
44633.6 19
0
10 2-In NAND~
219 656 1263 0 3 22
0 30 29 27
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U17A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
4299 0 0
2
44633.6 20
0
10 2-In NAND~
219 656 1168 0 3 22
0 29 32 28
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U17B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
9672 0 0
2
44633.6 21
0
9 Inverter~
13 432 1306 0 2 22
0 2 29
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U6B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 15 0
1 U
7876 0 0
2
44633.6 22
0
14 Logic Display~
6 890 1226 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
44633.6 23
0
14 Logic Display~
6 890 1659 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
44633.6 24
0
9 Inverter~
13 432 1739 0 2 22
0 2 11
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U6C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 15 0
1 U
7100 0 0
2
44633.6 25
0
10 2-In NAND~
219 656 1601 0 3 22
0 11 14 10
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U17C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
3820 0 0
2
44633.6 26
0
10 2-In NAND~
219 656 1696 0 3 22
0 12 11 9
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U17D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
7678 0 0
2
44633.6 27
0
10 2-In NAND~
219 800 1687 0 3 22
0 4 9 8
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
961 0 0
2
44633.6 28
0
10 2-In NAND~
219 800 1610 0 3 22
0 10 8 4
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 18 0
1 U
3178 0 0
2
44633.6 29
0
10 2-In NAND~
219 509 1610 0 3 22
0 15 12 14
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U18C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 18 0
1 U
3409 0 0
2
44633.6 30
0
10 2-In NAND~
219 510 1687 0 3 22
0 14 13 12
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U18D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 18 0
1 U
3951 0 0
2
44633.6 31
0
10 2-In NAND~
219 367 1696 0 3 22
0 2 16 13
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 19 0
1 U
8885 0 0
2
44633.6 32
0
10 2-In NAND~
219 368 1601 0 3 22
0 5 2 15
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 19 0
1 U
3780 0 0
2
44633.6 33
0
9 Inverter~
13 279 1642 0 2 22
0 5 16
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U6D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 15 0
1 U
9265 0 0
2
44633.6 34
0
9 Inverter~
13 279 1431 0 2 22
0 6 25
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 15 0
1 U
9442 0 0
2
44633.6 35
0
10 2-In NAND~
219 368 1390 0 3 22
0 6 2 24
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
9424 0 0
2
44633.6 36
0
10 2-In NAND~
219 367 1485 0 3 22
0 2 25 22
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U19D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
9968 0 0
2
44633.6 37
0
10 2-In NAND~
219 510 1476 0 3 22
0 23 22 21
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U20A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
9281 0 0
2
44633.6 38
0
10 2-In NAND~
219 509 1399 0 3 22
0 24 21 23
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U20B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 20 0
1 U
8464 0 0
2
44633.6 39
0
10 2-In NAND~
219 800 1399 0 3 22
0 19 17 5
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U20C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 20 0
1 U
7168 0 0
2
44633.6 40
0
10 2-In NAND~
219 800 1476 0 3 22
0 5 18 17
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U20D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 20 0
1 U
3171 0 0
2
44633.6 41
0
10 2-In NAND~
219 656 1485 0 3 22
0 21 20 18
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U21A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
4139 0 0
2
44633.6 42
0
10 2-In NAND~
219 656 1390 0 3 22
0 20 23 19
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U21B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
6435 0 0
2
44633.6 43
0
9 Inverter~
13 432 1528 0 2 22
0 2 20
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U6F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 15 0
1 U
5283 0 0
2
44633.6 44
0
14 Logic Display~
6 890 1448 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
44633.6 45
0
14 Logic Display~
6 1233 98 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
44633.6 46
0
14 Logic Display~
6 1282 98 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
44633.6 47
0
14 Logic Display~
6 1380 97 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
969 0 0
2
44633.6 48
0
14 Logic Display~
6 1331 97 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-8 -21 6 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8402 0 0
2
44633.6 49
0
14 Logic Display~
6 888 178 0 1 2
10 74
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3751 0 0
2
44633.6 50
0
9 Inverter~
13 430 258 0 2 22
0 2 77
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
4292 0 0
2
44633.6 51
0
10 2-In NAND~
219 654 120 0 3 22
0 77 80 76
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
6118 0 0
2
44633.6 52
0
10 2-In NAND~
219 654 215 0 3 22
0 78 77 75
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
34 0 0
2
44633.6 53
0
10 2-In NAND~
219 798 206 0 3 22
0 46 75 74
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
6357 0 0
2
44633.6 54
0
10 2-In NAND~
219 798 129 0 3 22
0 76 74 46
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
319 0 0
2
44633.6 55
0
10 2-In NAND~
219 507 129 0 3 22
0 81 78 80
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3976 0 0
2
44633.6 56
0
10 2-In NAND~
219 508 206 0 3 22
0 80 79 78
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7634 0 0
2
44633.6 57
0
10 2-In NAND~
219 365 215 0 3 22
0 2 82 79
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
523 0 0
2
44633.6 58
0
10 2-In NAND~
219 366 120 0 3 22
0 83 2 81
0
0 0 608 0
4 7400
-7 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
6748 0 0
2
44633.6 59
0
9 Inverter~
13 277 161 0 2 22
0 83 82
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6901 0 0
2
44633.6 60
0
9 Inverter~
13 277 372 0 2 22
0 46 73
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 U1E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
842 0 0
2
44633.6 61
0
10 2-In NAND~
219 366 331 0 3 22
0 46 2 72
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
3277 0 0
2
44633.6 62
0
10 2-In NAND~
219 365 426 0 3 22
0 2 73 70
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
4212 0 0
2
44633.6 63
0
10 2-In NAND~
219 508 417 0 3 22
0 71 70 69
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U10C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
4720 0 0
2
44633.6 64
0
10 2-In NAND~
219 507 340 0 3 22
0 72 69 71
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U10D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
5551 0 0
2
44633.6 65
0
10 2-In NAND~
219 798 340 0 3 22
0 67 65 45
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
6986 0 0
2
44633.6 66
0
10 2-In NAND~
219 798 417 0 3 22
0 45 66 65
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U11B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
8745 0 0
2
44633.6 67
0
10 2-In NAND~
219 654 426 0 3 22
0 69 68 66
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U11C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
9592 0 0
2
44633.6 68
0
10 2-In NAND~
219 654 331 0 3 22
0 68 71 67
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U11D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
8748 0 0
2
44633.6 69
0
9 Inverter~
13 430 469 0 2 22
0 2 68
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
7168 0 0
2
44633.6 70
0
14 Logic Display~
6 888 389 0 1 2
10 65
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
631 0 0
2
44633.6 71
0
14 Logic Display~
6 888 822 0 1 2
10 47
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9466 0 0
2
44633.6 72
0
9 Inverter~
13 430 902 0 2 22
0 2 50
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U12A
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
3266 0 0
2
44633.6 73
0
10 2-In NAND~
219 654 764 0 3 22
0 50 53 49
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
7693 0 0
2
44633.6 74
0
10 2-In NAND~
219 654 859 0 3 22
0 51 50 48
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
3723 0 0
2
44633.6 75
0
10 2-In NAND~
219 798 850 0 3 22
0 3 48 47
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U13C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3440 0 0
2
44633.6 76
0
10 2-In NAND~
219 798 773 0 3 22
0 49 47 3
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U13D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
6263 0 0
2
44633.6 77
0
10 2-In NAND~
219 507 773 0 3 22
0 54 51 53
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
4900 0 0
2
44633.6 78
0
10 2-In NAND~
219 508 850 0 3 22
0 53 52 51
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
8783 0 0
2
44633.6 79
0
10 2-In NAND~
219 365 859 0 3 22
0 2 55 52
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3221 0 0
2
44633.6 80
0
10 2-In NAND~
219 366 764 0 3 22
0 44 2 54
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
3215 0 0
2
44633.6 81
0
9 Inverter~
13 277 805 0 2 22
0 44 55
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U12B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
7903 0 0
2
44633.6 82
0
9 Inverter~
13 277 594 0 2 22
0 45 64
0
0 0 608 270
6 74LS04
-21 -19 21 -11
4 U12C
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
7121 0 0
2
44633.6 83
0
10 2-In NAND~
219 366 553 0 3 22
0 45 2 63
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
4484 0 0
2
44633.6 84
0
10 2-In NAND~
219 365 648 0 3 22
0 2 64 61
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
5996 0 0
2
44633.6 85
0
10 2-In NAND~
219 508 639 0 3 22
0 62 61 60
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U15C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
7804 0 0
2
44633.6 86
0
10 2-In NAND~
219 507 562 0 3 22
0 63 60 62
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U15D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
5523 0 0
2
44633.6 87
0
10 2-In NAND~
219 798 562 0 3 22
0 58 56 44
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
3330 0 0
2
44633.6 88
0
10 2-In NAND~
219 798 639 0 3 22
0 44 57 56
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
3465 0 0
2
44633.6 89
0
10 2-In NAND~
219 654 648 0 3 22
0 60 59 57
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
8396 0 0
2
44633.6 90
0
10 2-In NAND~
219 654 553 0 3 22
0 59 62 58
0
0 0 608 0
4 7400
-7 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
3685 0 0
2
44633.6 91
0
9 Inverter~
13 430 691 0 2 22
0 2 59
0
0 0 608 0
6 74LS04
-21 -19 21 -11
4 U12D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
7849 0 0
2
44633.6 92
0
14 Logic Display~
6 888 611 0 1 2
10 56
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6343 0 0
2
44633.6 93
0
14 Logic Display~
6 1021 100 0 1 2
10 46
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
44633.6 94
0
14 Logic Display~
6 1074 100 0 1 2
10 45
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
44633.6 95
0
14 Logic Display~
6 1181 100 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5776 0 0
2
44633.6 96
0
14 Logic Display~
6 1127 101 0 1 2
10 44
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7207 0 0
2
44633.6 97
0
160
0 0 2 0 0 8192 0 0 0 26 10 3
327 1739
142 1739
142 1528
1 0 3 0 0 4096 0 12 0 0 80 4
344 948
287 948
287 949
282 949
1 0 4 0 0 4224 0 49 0 0 13 3
1380 115
1380 1610
859 1610
1 0 5 0 0 4224 0 50 0 0 7 3
1331 115
1331 1399
923 1399
1 0 6 0 0 4224 0 48 0 0 8 3
1282 116
1282 1177
923 1177
1 0 7 0 0 4224 0 47 0 0 9 3
1233 116
1233 966
923 966
0 0 5 0 0 0 0 0 0 30 29 5
859 1399
923 1399
923 1561
282 1561
282 1592
0 0 6 0 0 0 0 0 0 47 46 5
859 1177
923 1177
923 1345
282 1345
282 1381
0 0 7 0 0 0 0 0 0 64 63 5
859 966
923 966
923 1126
282 1126
282 1159
0 0 2 0 0 8192 0 0 0 43 11 3
327 1528
142 1528
142 1306
0 0 2 0 0 0 0 0 0 60 12 3
327 1306
142 1306
142 1095
0 0 2 0 0 0 0 0 0 77 81 3
327 1095
142 1095
142 901
1 3 4 0 0 0 0 29 30 0 0 6
776 1678
767 1678
767 1653
859 1653
859 1610
827 1610
2 0 8 0 0 12416 0 30 0 0 15 5
776 1619
767 1619
767 1643
846 1643
846 1687
3 1 8 0 0 0 0 29 25 0 0 3
827 1687
890 1687
890 1677
3 2 9 0 0 4224 0 28 29 0 0 2
683 1696
776 1696
3 1 10 0 0 4224 0 27 30 0 0 2
683 1601
776 1601
2 0 11 0 0 4096 0 28 0 0 23 2
632 1705
607 1705
2 0 12 0 0 12288 0 31 0 0 20 5
485 1619
476 1619
476 1643
555 1643
555 1687
3 1 12 0 0 4224 0 32 28 0 0 2
537 1687
632 1687
3 2 13 0 0 4224 0 33 32 0 0 2
394 1696
486 1696
1 0 14 0 0 12288 0 32 0 0 24 5
486 1678
476 1678
476 1653
568 1653
568 1610
2 1 11 0 0 4224 0 26 27 0 0 4
453 1739
607 1739
607 1592
632 1592
3 2 14 0 0 4224 0 31 27 0 0 2
536 1610
632 1610
3 1 15 0 0 4224 0 34 31 0 0 2
395 1601
485 1601
1 0 2 0 0 0 0 26 0 0 27 3
417 1739
327 1739
327 1687
1 2 2 0 0 0 0 33 34 0 0 4
343 1687
327 1687
327 1610
344 1610
2 2 16 0 0 8320 0 35 33 0 0 3
282 1660
282 1705
343 1705
1 1 5 0 0 0 0 35 34 0 0 3
282 1624
282 1592
344 1592
1 3 5 0 0 0 0 42 41 0 0 6
776 1467
767 1467
767 1442
859 1442
859 1399
827 1399
2 0 17 0 0 12416 0 41 0 0 32 5
776 1408
767 1408
767 1432
846 1432
846 1476
3 1 17 0 0 0 0 42 46 0 0 3
827 1476
890 1476
890 1466
3 2 18 0 0 4224 0 43 42 0 0 2
683 1485
776 1485
3 1 19 0 0 4224 0 44 41 0 0 2
683 1390
776 1390
2 0 20 0 0 4096 0 43 0 0 40 2
632 1494
607 1494
2 0 21 0 0 12288 0 40 0 0 37 5
485 1408
476 1408
476 1432
555 1432
555 1476
3 1 21 0 0 4224 0 39 43 0 0 2
537 1476
632 1476
3 2 22 0 0 4224 0 38 39 0 0 2
394 1485
486 1485
1 0 23 0 0 12288 0 39 0 0 41 5
486 1467
476 1467
476 1442
568 1442
568 1399
2 1 20 0 0 4224 0 45 44 0 0 4
453 1528
607 1528
607 1381
632 1381
3 2 23 0 0 4224 0 40 44 0 0 2
536 1399
632 1399
3 1 24 0 0 4224 0 37 40 0 0 2
395 1390
485 1390
1 0 2 0 0 0 0 45 0 0 44 3
417 1528
327 1528
327 1476
1 2 2 0 0 0 0 38 37 0 0 4
343 1476
327 1476
327 1399
344 1399
2 2 25 0 0 8320 0 36 38 0 0 3
282 1449
282 1494
343 1494
1 1 6 0 0 0 0 36 37 0 0 3
282 1413
282 1381
344 1381
1 3 6 0 0 0 0 20 19 0 0 6
776 1245
767 1245
767 1220
859 1220
859 1177
827 1177
2 0 26 0 0 12416 0 19 0 0 49 5
776 1186
767 1186
767 1210
846 1210
846 1254
3 1 26 0 0 0 0 20 24 0 0 3
827 1254
890 1254
890 1244
3 2 27 0 0 4224 0 21 20 0 0 2
683 1263
776 1263
3 1 28 0 0 4224 0 22 19 0 0 2
683 1168
776 1168
2 0 29 0 0 4096 0 21 0 0 57 2
632 1272
607 1272
2 0 30 0 0 12288 0 18 0 0 54 5
485 1186
476 1186
476 1210
555 1210
555 1254
3 1 30 0 0 4224 0 17 21 0 0 2
537 1254
632 1254
3 2 31 0 0 4224 0 16 17 0 0 2
394 1263
486 1263
1 0 32 0 0 12288 0 17 0 0 58 5
486 1245
476 1245
476 1220
568 1220
568 1177
2 1 29 0 0 4224 0 23 22 0 0 4
453 1306
607 1306
607 1159
632 1159
3 2 32 0 0 4224 0 18 22 0 0 2
536 1177
632 1177
3 1 33 0 0 4224 0 15 18 0 0 2
395 1168
485 1168
1 0 2 0 0 0 0 23 0 0 61 3
417 1306
327 1306
327 1254
1 2 2 0 0 0 0 16 15 0 0 4
343 1254
327 1254
327 1177
344 1177
2 2 34 0 0 8320 0 14 16 0 0 3
282 1227
282 1272
343 1272
1 1 7 0 0 0 0 14 15 0 0 3
282 1191
282 1159
344 1159
1 3 7 0 0 0 0 7 8 0 0 6
776 1034
767 1034
767 1009
859 1009
859 966
827 966
2 0 35 0 0 12416 0 8 0 0 66 5
776 975
767 975
767 999
846 999
846 1043
3 1 35 0 0 0 0 7 3 0 0 3
827 1043
890 1043
890 1033
3 2 36 0 0 4224 0 6 7 0 0 2
683 1052
776 1052
3 1 37 0 0 4224 0 5 8 0 0 2
683 957
776 957
2 0 38 0 0 4096 0 6 0 0 74 2
632 1061
607 1061
2 0 39 0 0 12288 0 9 0 0 71 5
485 975
476 975
476 999
555 999
555 1043
3 1 39 0 0 4224 0 10 6 0 0 2
537 1043
632 1043
3 2 40 0 0 4224 0 11 10 0 0 2
394 1052
486 1052
1 0 41 0 0 12288 0 10 0 0 75 5
486 1034
476 1034
476 1009
568 1009
568 966
2 1 38 0 0 4224 0 4 5 0 0 4
453 1095
607 1095
607 948
632 948
3 2 41 0 0 4224 0 9 5 0 0 2
536 966
632 966
3 1 42 0 0 4224 0 12 9 0 0 2
395 957
485 957
1 0 2 0 0 0 0 4 0 0 78 3
417 1095
327 1095
327 1043
1 2 2 0 0 0 0 11 12 0 0 4
343 1043
327 1043
327 966
344 966
2 2 43 0 0 8320 0 13 11 0 0 3
282 1016
282 1061
343 1061
1 0 3 0 0 16384 0 13 0 0 82 6
282 980
282 948
281 948
281 923
924 923
924 773
1 0 2 0 0 8320 0 1 0 0 105 5
93 111
142 111
142 901
325 901
325 902
1 0 3 0 0 4224 0 97 0 0 92 3
1181 118
1181 773
857 773
1 0 44 0 0 4096 0 98 0 0 86 3
1127 119
1127 562
921 562
1 0 45 0 0 4096 0 96 0 0 87 3
1074 118
1074 340
921 340
1 0 46 0 0 8192 0 95 0 0 88 3
1021 118
1021 129
921 129
0 0 44 0 0 12416 0 0 0 109 108 5
857 562
921 562
921 724
280 724
280 755
0 0 45 0 0 12416 0 0 0 126 125 5
857 340
921 340
921 508
280 508
280 544
0 0 46 0 0 12416 0 0 0 143 142 5
857 129
921 129
921 289
280 289
280 322
0 0 2 0 0 0 0 0 0 122 81 2
325 691
142 691
0 0 2 0 0 0 0 0 0 139 81 2
325 469
142 469
0 0 2 0 0 0 0 0 0 156 81 2
325 258
142 258
1 3 3 0 0 0 0 77 78 0 0 6
774 841
765 841
765 816
857 816
857 773
825 773
2 0 47 0 0 12416 0 78 0 0 94 5
774 782
765 782
765 806
844 806
844 850
3 1 47 0 0 0 0 77 73 0 0 3
825 850
888 850
888 840
3 2 48 0 0 4224 0 76 77 0 0 2
681 859
774 859
3 1 49 0 0 4224 0 75 78 0 0 2
681 764
774 764
2 0 50 0 0 4096 0 76 0 0 102 2
630 868
605 868
2 0 51 0 0 12288 0 79 0 0 99 5
483 782
474 782
474 806
553 806
553 850
3 1 51 0 0 4224 0 80 76 0 0 2
535 850
630 850
3 2 52 0 0 4224 0 81 80 0 0 2
392 859
484 859
1 0 53 0 0 12288 0 80 0 0 103 5
484 841
474 841
474 816
566 816
566 773
2 1 50 0 0 4224 0 74 75 0 0 4
451 902
605 902
605 755
630 755
3 2 53 0 0 4224 0 79 75 0 0 2
534 773
630 773
3 1 54 0 0 4224 0 82 79 0 0 2
393 764
483 764
1 0 2 0 0 0 0 74 0 0 106 3
415 902
325 902
325 850
1 2 2 0 0 0 0 81 82 0 0 4
341 850
325 850
325 773
342 773
2 2 55 0 0 8320 0 83 81 0 0 3
280 823
280 868
341 868
1 1 44 0 0 0 0 83 82 0 0 3
280 787
280 755
342 755
1 3 44 0 0 0 0 90 89 0 0 6
774 630
765 630
765 605
857 605
857 562
825 562
2 0 56 0 0 12416 0 89 0 0 111 5
774 571
765 571
765 595
844 595
844 639
3 1 56 0 0 0 0 90 94 0 0 3
825 639
888 639
888 629
3 2 57 0 0 4224 0 91 90 0 0 2
681 648
774 648
3 1 58 0 0 4224 0 92 89 0 0 2
681 553
774 553
2 0 59 0 0 4096 0 91 0 0 119 2
630 657
605 657
2 0 60 0 0 12288 0 88 0 0 116 5
483 571
474 571
474 595
553 595
553 639
3 1 60 0 0 4224 0 87 91 0 0 2
535 639
630 639
3 2 61 0 0 4224 0 86 87 0 0 2
392 648
484 648
1 0 62 0 0 12288 0 87 0 0 120 5
484 630
474 630
474 605
566 605
566 562
2 1 59 0 0 4224 0 93 92 0 0 4
451 691
605 691
605 544
630 544
3 2 62 0 0 4224 0 88 92 0 0 2
534 562
630 562
3 1 63 0 0 4224 0 85 88 0 0 2
393 553
483 553
1 0 2 0 0 0 0 93 0 0 123 3
415 691
325 691
325 639
1 2 2 0 0 0 0 86 85 0 0 4
341 639
325 639
325 562
342 562
2 2 64 0 0 8320 0 84 86 0 0 3
280 612
280 657
341 657
1 1 45 0 0 0 0 84 85 0 0 3
280 576
280 544
342 544
1 3 45 0 0 0 0 68 67 0 0 6
774 408
765 408
765 383
857 383
857 340
825 340
2 0 65 0 0 12416 0 67 0 0 128 5
774 349
765 349
765 373
844 373
844 417
3 1 65 0 0 0 0 68 72 0 0 3
825 417
888 417
888 407
3 2 66 0 0 4224 0 69 68 0 0 2
681 426
774 426
3 1 67 0 0 4224 0 70 67 0 0 2
681 331
774 331
2 0 68 0 0 4096 0 69 0 0 136 2
630 435
605 435
2 0 69 0 0 12288 0 66 0 0 133 5
483 349
474 349
474 373
553 373
553 417
3 1 69 0 0 4224 0 65 69 0 0 2
535 417
630 417
3 2 70 0 0 4224 0 64 65 0 0 2
392 426
484 426
1 0 71 0 0 12288 0 65 0 0 137 5
484 408
474 408
474 383
566 383
566 340
2 1 68 0 0 4224 0 71 70 0 0 4
451 469
605 469
605 322
630 322
3 2 71 0 0 4224 0 66 70 0 0 2
534 340
630 340
3 1 72 0 0 4224 0 63 66 0 0 2
393 331
483 331
1 0 2 0 0 0 0 71 0 0 140 3
415 469
325 469
325 417
1 2 2 0 0 0 0 64 63 0 0 4
341 417
325 417
325 340
342 340
2 2 73 0 0 8320 0 62 64 0 0 3
280 390
280 435
341 435
1 1 46 0 0 0 0 62 63 0 0 3
280 354
280 322
342 322
1 3 46 0 0 0 0 55 56 0 0 6
774 197
765 197
765 172
857 172
857 129
825 129
2 0 74 0 0 12416 0 56 0 0 145 5
774 138
765 138
765 162
844 162
844 206
3 1 74 0 0 0 0 55 51 0 0 3
825 206
888 206
888 196
3 2 75 0 0 4224 0 54 55 0 0 2
681 215
774 215
3 1 76 0 0 4224 0 53 56 0 0 2
681 120
774 120
2 0 77 0 0 4096 0 54 0 0 153 2
630 224
605 224
2 0 78 0 0 12288 0 57 0 0 150 5
483 138
474 138
474 162
553 162
553 206
3 1 78 0 0 4224 0 58 54 0 0 2
535 206
630 206
3 2 79 0 0 4224 0 59 58 0 0 2
392 215
484 215
1 0 80 0 0 12288 0 58 0 0 154 5
484 197
474 197
474 172
566 172
566 129
2 1 77 0 0 4224 0 52 53 0 0 4
451 258
605 258
605 111
630 111
3 2 80 0 0 4224 0 57 53 0 0 2
534 129
630 129
3 1 81 0 0 4224 0 60 57 0 0 2
393 120
483 120
1 0 2 0 0 0 0 52 0 0 157 3
415 258
325 258
325 206
1 2 2 0 0 0 0 59 60 0 0 4
341 206
325 206
325 129
342 129
2 2 82 0 0 8320 0 61 59 0 0 3
280 179
280 224
341 224
1 0 83 0 0 4096 0 61 0 0 160 2
280 143
280 111
1 1 83 0 0 4224 0 2 60 0 0 2
218 111
342 111
42
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1362 39 1394 63
1371 48 1384 64
2 Q8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1314 40 1346 64
1323 49 1336 65
2 Q7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1264 42 1296 66
1273 51 1286 67
2 Q6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1216 41 1248 65
1225 50 1238 66
2 Q5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
694 1633 755 1657
704 1641 744 1657
5 SLAVE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
690 1422 751 1446
700 1430 740 1446
5 SLAVE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
397 1635 466 1659
407 1643 455 1659
6 MASTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
393 1424 462 1448
403 1432 451 1448
6 MASTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
693 1199 754 1223
703 1207 743 1223
5 SLAVE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
689 988 750 1012
699 996 739 1012
5 SLAVE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
396 1201 465 1225
406 1209 454 1225
6 MASTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
392 990 461 1014
402 998 450 1014
6 MASTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
895 1646 926 1668
902 1653 918 1669
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
896 1580 919 1602
903 1587 911 1603
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
896 1370 919 1392
903 1377 911 1393
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
895 1436 926 1458
902 1443 918 1459
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
896 1149 919 1171
903 1156 911 1172
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
895 1215 926 1237
902 1222 918 1238
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
895 1005 926 1027
902 1012 918 1028
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
896 939 919 961
903 946 911 962
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
692 796 753 820
702 804 742 820
5 SLAVE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
688 585 749 609
698 593 738 609
5 SLAVE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
395 798 464 822
405 806 453 822
6 MASTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
391 587 460 611
401 595 449 611
6 MASTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
691 362 752 386
701 370 741 386
5 SLAVE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
687 151 748 175
697 159 737 175
5 SLAVE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
394 364 463 388
404 372 452 388
6 MASTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
390 153 459 177
400 161 448 177
6 MASTER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
893 809 924 831
900 816 916 832
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
894 743 917 765
901 750 909 766
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
894 533 917 555
901 540 909 556
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
893 599 924 621
900 606 916 622
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
894 312 917 334
901 319 909 335
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
893 378 924 400
900 385 916 401
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
893 168 924 190
900 175 916 191
2 Q'
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
894 102 917 124
901 109 909 125
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1165 43 1198 65
1173 50 1189 66
2 Q4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1112 43 1143 65
1119 50 1135 66
2 Q3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1057 43 1090 65
1065 50 1081 66
2 Q2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1005 41 1036 63
1012 49 1028 65
2 Q1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1145 18 1260 40
1154 25 1250 41
12 PARALLEL OUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 23
53 26 247 49
63 36 236 51
23 RANGKAIAN REGISTER SIPO
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
